magic
tech sky130A
magscale 1 2
timestamp 1729239461
<< pwell >>
rect -196 -503 1126 491
<< psubdiff >>
rect -176 436 -116 470
rect 1046 436 1106 470
rect -176 410 -142 436
rect 1072 410 1106 436
rect -176 -449 -142 -423
rect 1072 -449 1106 -423
rect -176 -483 -116 -449
rect 1046 -483 1106 -449
<< psubdiffcont >>
rect -116 436 1046 470
rect -176 -423 -142 410
rect 1072 -423 1106 410
rect -116 -483 1046 -449
<< poly >>
rect -92 389 0 405
rect -92 355 -76 389
rect -42 355 0 389
rect -92 339 0 355
rect -30 296 0 339
rect 930 386 1022 402
rect 930 352 972 386
rect 1006 352 1022 386
rect 930 336 1022 352
rect 930 302 960 336
rect 58 -42 872 1
rect -30 -352 0 -345
rect -92 -368 0 -352
rect -92 -402 -76 -368
rect -42 -402 0 -368
rect -92 -418 0 -402
rect 930 -352 960 -332
rect 930 -368 1022 -352
rect 930 -402 972 -368
rect 1006 -402 1022 -368
rect 930 -418 1022 -402
<< polycont >>
rect -76 355 -42 389
rect 972 352 1006 386
rect -76 -402 -42 -368
rect 972 -402 1006 -368
<< locali >>
rect -176 436 -116 470
rect 1046 436 1106 470
rect -176 410 -142 436
rect 1072 410 1106 436
rect -92 355 -76 389
rect -42 355 -26 389
rect -76 276 -42 355
rect 956 352 972 386
rect 1006 352 1022 386
rect 972 276 1006 352
rect -76 -368 -42 -318
rect 972 -368 1006 -318
rect -92 -402 -76 -368
rect -42 -402 -26 -368
rect 956 -402 972 -368
rect 1006 -402 1022 -368
rect -176 -449 -142 -423
rect 1072 -449 1106 -423
rect -176 -483 -116 -449
rect 1046 -483 1106 -449
<< viali >>
rect 230 436 264 470
rect 665 436 699 470
rect -76 355 -42 389
rect 972 352 1006 386
rect -76 -402 -42 -368
rect 972 -402 1006 -368
rect 230 -483 264 -449
rect 666 -483 700 -449
<< metal1 >>
rect 208 424 218 484
rect 276 424 286 484
rect 643 423 653 483
rect 711 423 721 483
rect -88 389 -30 395
rect -88 355 -76 389
rect -42 355 -30 389
rect -88 349 -30 355
rect 960 386 1018 392
rect 960 352 972 386
rect 1006 352 1018 386
rect -82 289 -36 349
rect 960 346 1018 352
rect -82 88 52 289
rect 208 88 218 289
rect 276 88 286 289
rect 426 88 436 290
rect 494 88 504 290
rect 6 56 52 88
rect 645 87 655 289
rect 711 87 721 289
rect 967 288 1012 346
rect 878 88 1012 288
rect 878 56 924 88
rect 6 10 138 56
rect 792 10 924 56
rect 356 -98 574 -52
rect -82 -130 53 -129
rect -82 -330 0 -130
rect 58 -330 68 -130
rect -82 -362 -36 -330
rect 208 -331 218 -130
rect 276 -331 286 -130
rect 442 -330 488 -98
rect 878 -130 1013 -129
rect 644 -331 654 -130
rect 712 -331 722 -130
rect 862 -330 872 -130
rect 930 -330 1013 -130
rect 966 -362 1012 -330
rect -88 -368 -30 -362
rect -88 -402 -76 -368
rect -42 -402 -30 -368
rect -88 -408 -30 -402
rect 960 -368 1018 -362
rect 960 -402 972 -368
rect 1006 -402 1018 -368
rect 960 -408 1018 -402
rect 208 -496 218 -436
rect 276 -496 286 -436
rect 644 -496 654 -436
rect 712 -496 722 -436
<< via1 >>
rect 218 470 276 484
rect 218 436 230 470
rect 230 436 264 470
rect 264 436 276 470
rect 218 424 276 436
rect 653 470 711 483
rect 653 436 665 470
rect 665 436 699 470
rect 699 436 711 470
rect 653 423 711 436
rect 218 88 276 289
rect 436 88 494 290
rect 655 87 711 289
rect 0 -330 58 -130
rect 218 -331 276 -130
rect 654 -331 712 -130
rect 872 -330 930 -130
rect 218 -449 276 -436
rect 218 -483 230 -449
rect 230 -483 264 -449
rect 264 -483 276 -449
rect 218 -496 276 -483
rect 654 -449 712 -436
rect 654 -483 666 -449
rect 666 -483 700 -449
rect 700 -483 712 -449
rect 654 -496 712 -483
<< metal2 >>
rect 218 484 276 494
rect 218 414 276 424
rect 653 483 711 493
rect 227 329 267 414
rect 653 413 711 423
rect 657 341 709 413
rect 218 289 276 329
rect 218 78 276 88
rect 436 290 494 300
rect 436 49 494 88
rect 655 289 711 341
rect 655 77 711 87
rect 446 -3 485 49
rect 10 -42 920 -3
rect 10 -120 49 -42
rect 881 -120 920 -42
rect 0 -130 58 -120
rect 0 -340 58 -330
rect 218 -130 276 -120
rect 218 -372 276 -331
rect 654 -130 712 -120
rect 227 -426 268 -372
rect 654 -373 712 -331
rect 872 -130 930 -120
rect 872 -340 930 -330
rect 662 -426 704 -373
rect 218 -436 276 -426
rect 218 -506 276 -496
rect 654 -436 712 -426
rect 654 -506 712 -496
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729239461
transform 1 0 -15 0 1 -230
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729239461
transform 1 0 -15 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729239461
transform 1 0 945 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_4
timestamp 1729239461
transform 1 0 945 0 1 -230
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_HRGC9X  sky130_fd_pr__nfet_01v8_HRGC9X_0
timestamp 1729239461
transform 1 0 465 0 1 -230
box -465 -188 465 188
use sky130_fd_pr__nfet_01v8_HRGC9X  sky130_fd_pr__nfet_01v8_HRGC9X_1
timestamp 1729239461
transform 1 0 465 0 1 188
box -465 -188 465 188
<< labels >>
flabel metal1 29 35 29 35 0 FreeSans 160 0 0 0 D8
port 0 nsew
flabel psubdiffcont -53 -467 -53 -467 0 FreeSans 160 0 0 0 GND
port 1 nsew
flabel metal2 31 -78 31 -78 0 FreeSans 160 0 0 0 OUT
port 2 nsew
<< end >>
