magic
tech sky130A
magscale 1 2
timestamp 1729169387
<< nwell >>
rect -176 53 822 1391
rect -176 19 306 53
rect 599 19 822 53
rect -176 -1489 822 19
<< nsubdiff >>
rect -140 1321 -80 1355
rect 726 1321 786 1355
rect -140 1295 -106 1321
rect 752 1295 786 1321
rect -140 -1419 -106 -1393
rect 752 -1419 786 -1393
rect -140 -1453 -80 -1419
rect 726 -1453 786 -1419
<< nsubdiffcont >>
rect -80 1321 726 1355
rect -140 -1393 -106 1295
rect 752 -1393 786 1295
rect -80 -1453 726 -1419
<< poly >>
rect -56 1282 36 1298
rect -56 1248 -40 1282
rect -6 1248 36 1282
rect -56 1232 36 1248
rect 6 1211 36 1232
rect 610 1283 702 1299
rect 610 1249 652 1283
rect 686 1249 702 1283
rect 610 1233 702 1249
rect 610 1212 640 1233
rect 94 597 294 703
rect -56 581 36 597
rect -56 547 -40 581
rect -6 547 36 581
rect -56 531 36 547
rect 6 510 36 531
rect 610 581 702 597
rect 610 547 652 581
rect 686 547 702 581
rect 610 531 702 547
rect 610 510 640 531
rect 94 -103 552 3
rect 6 -631 36 -610
rect -56 -647 36 -631
rect -56 -681 -40 -647
rect -6 -681 36 -647
rect -56 -697 36 -681
rect 610 -631 640 -610
rect 610 -647 702 -631
rect 610 -681 652 -647
rect 686 -681 702 -647
rect 610 -697 702 -681
rect 353 -803 553 -697
rect 6 -1331 36 -1310
rect -56 -1347 36 -1331
rect -56 -1381 -40 -1347
rect -6 -1381 36 -1347
rect -56 -1397 36 -1381
rect 610 -1331 640 -1310
rect 610 -1347 702 -1331
rect 610 -1381 652 -1347
rect 686 -1381 702 -1347
rect 610 -1397 702 -1381
<< polycont >>
rect -40 1248 -6 1282
rect 652 1249 686 1283
rect -40 547 -6 581
rect 652 547 686 581
rect -40 -681 -6 -647
rect 652 -681 686 -647
rect -40 -1381 -6 -1347
rect 652 -1381 686 -1347
<< locali >>
rect -140 1321 -80 1355
rect 726 1321 786 1355
rect -140 1295 -106 1321
rect 752 1295 786 1321
rect -56 1248 -40 1282
rect -6 1248 10 1282
rect 636 1249 652 1283
rect 686 1249 702 1283
rect -56 547 -40 581
rect -6 547 10 581
rect 636 547 652 581
rect 686 547 702 581
rect -56 -681 -40 -647
rect -6 -681 10 -647
rect 636 -681 652 -647
rect 686 -681 702 -647
rect -56 -1381 -40 -1347
rect -6 -1381 10 -1347
rect 636 -1381 652 -1347
rect 686 -1381 702 -1347
rect -140 -1419 -106 -1393
rect 752 -1419 786 -1393
rect -140 -1453 -80 -1419
rect 726 -1453 786 -1419
<< viali >>
rect 652 1321 686 1355
rect -40 1248 -6 1282
rect 652 1249 686 1283
rect -40 547 -6 581
rect 652 547 686 581
rect -40 -681 -6 -647
rect 652 -681 686 -647
rect -40 -1381 -6 -1347
rect 652 -1381 686 -1347
rect -40 -1453 -6 -1419
<< metal1 >>
rect 640 1355 698 1361
rect 640 1321 652 1355
rect 686 1321 698 1355
rect -52 1282 6 1288
rect -52 1248 -40 1282
rect -6 1248 6 1282
rect -52 1242 6 1248
rect 640 1283 698 1321
rect 640 1249 652 1283
rect 686 1249 698 1283
rect 640 1243 698 1249
rect -40 1200 -6 1242
rect 652 1200 686 1243
rect -46 1188 88 1200
rect -59 812 -49 1188
rect 3 812 88 1188
rect -46 800 88 812
rect 306 754 340 848
rect 558 800 692 1200
rect 563 754 598 800
rect 306 719 598 754
rect -52 581 6 587
rect -52 547 -40 581
rect -6 547 6 581
rect -52 541 6 547
rect -40 500 -6 541
rect -46 488 88 500
rect -46 112 39 488
rect 91 112 101 488
rect -46 100 88 112
rect 47 -154 168 -119
rect 47 -200 82 -154
rect -45 -600 89 -200
rect -40 -641 -6 -600
rect -52 -647 6 -641
rect -52 -681 -40 -647
rect -6 -681 6 -647
rect -52 -687 6 -681
rect 306 -819 340 719
rect 640 581 698 587
rect 640 547 652 581
rect 686 547 698 581
rect 640 541 698 547
rect 652 500 686 541
rect 558 100 692 500
rect 564 54 599 100
rect 477 19 599 54
rect 558 -212 692 -200
rect 545 -588 555 -212
rect 607 -588 692 -212
rect 558 -600 692 -588
rect 652 -641 686 -600
rect 640 -647 698 -641
rect 640 -681 652 -647
rect 686 -681 698 -647
rect 640 -687 698 -681
rect 48 -853 340 -819
rect 48 -900 82 -853
rect -46 -1300 88 -900
rect 306 -948 340 -853
rect 558 -912 692 -900
rect 558 -1288 643 -912
rect 695 -1288 705 -912
rect 558 -1300 692 -1288
rect -40 -1341 -6 -1300
rect 652 -1341 686 -1300
rect -52 -1347 6 -1341
rect -52 -1381 -40 -1347
rect -6 -1381 6 -1347
rect -52 -1419 6 -1381
rect 640 -1347 698 -1341
rect 640 -1381 652 -1347
rect 686 -1381 698 -1347
rect 640 -1387 698 -1381
rect -52 -1453 -40 -1419
rect -6 -1453 6 -1419
rect -52 -1459 6 -1453
<< via1 >>
rect -49 812 3 1188
rect 39 112 91 488
rect 555 -588 607 -212
rect 643 -1288 695 -912
<< metal2 >>
rect -49 1188 3 1198
rect -53 812 -49 1188
rect 3 812 7 1188
rect -53 684 7 812
rect -53 628 -51 684
rect 5 628 7 684
rect -53 -726 7 628
rect 639 686 699 695
rect 639 617 699 626
rect 39 488 91 498
rect 39 102 91 112
rect 43 -16 86 102
rect 43 -84 602 -16
rect 559 -202 602 -84
rect 555 -212 607 -202
rect 555 -598 607 -588
rect 643 -728 695 617
rect 632 -784 641 -728
rect 697 -784 706 -728
rect -53 -795 7 -786
rect 643 -912 695 -784
rect 643 -1298 695 -1288
<< via2 >>
rect -51 628 5 684
rect 639 626 699 686
rect -53 -786 7 -726
rect 641 -784 697 -728
<< metal3 >>
rect -56 686 10 689
rect 634 686 704 691
rect -56 684 639 686
rect -56 628 -51 684
rect 5 628 639 684
rect -56 626 639 628
rect 699 626 704 686
rect -56 623 10 626
rect 634 621 704 626
rect -58 -726 12 -721
rect 636 -726 702 -723
rect -58 -786 -53 -726
rect 7 -728 702 -726
rect 7 -784 641 -728
rect 697 -784 702 -728
rect 7 -786 702 -784
rect -58 -791 12 -786
rect 636 -789 702 -786
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729158395
transform 1 0 21 0 1 -1100
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729158395
transform 1 0 21 0 1 1000
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729158395
transform 1 0 625 0 1 1000
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729158395
transform 1 0 625 0 1 300
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729158395
transform 1 0 21 0 1 300
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729158395
transform 1 0 21 0 1 -400
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729158395
transform 1 0 625 0 1 -400
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729158395
transform 1 0 625 0 1 -1100
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729158395
transform 1 0 323 0 1 1000
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729158395
transform 1 0 323 0 1 300
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729158395
transform 1 0 323 0 1 -400
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729158395
transform 1 0 323 0 1 -1100
box -323 -300 323 300
<< labels >>
flabel viali 668 1336 668 1336 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel metal1 586 74 586 74 0 FreeSans 160 0 0 0 D2
port 1 nsew
flabel metal2 62 22 62 22 0 FreeSans 160 0 0 0 D1
port 2 nsew
flabel viali -22 1266 -22 1266 0 FreeSans 160 0 0 0 D5
port 3 nsew
<< end >>
