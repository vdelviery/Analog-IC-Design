magic
tech sky130A
magscale 1 2
timestamp 1729402320
<< nwell >>
rect -176 -743 938 489
<< nsubdiff >>
rect -140 419 -80 453
rect 842 419 902 453
rect -140 393 -106 419
rect 868 393 902 419
rect -140 -673 -106 -647
rect 868 -673 902 -647
rect -140 -707 -80 -673
rect 842 -707 902 -673
<< nsubdiffcont >>
rect -80 419 842 453
rect -140 -647 -106 393
rect 868 -647 902 393
rect -80 -707 842 -673
<< poly >>
rect -56 381 36 397
rect -56 347 -40 381
rect -6 347 36 381
rect -56 331 36 347
rect 6 300 36 331
rect 726 381 818 397
rect 726 347 768 381
rect 802 347 818 381
rect 726 331 818 347
rect 726 300 756 331
rect 352 -323 410 -257
rect 6 -585 36 -554
rect -56 -601 36 -585
rect -56 -635 -40 -601
rect -6 -635 36 -601
rect -56 -651 36 -635
rect 726 -585 756 -554
rect 726 -601 818 -585
rect 726 -635 768 -601
rect 802 -635 818 -601
rect 726 -651 818 -635
<< polycont >>
rect -40 347 -6 381
rect 768 347 802 381
rect -40 -635 -6 -601
rect 768 -635 802 -601
<< locali >>
rect -140 419 -80 453
rect 842 419 902 453
rect -140 393 -106 419
rect 868 393 902 419
rect -56 347 -40 381
rect -6 347 10 381
rect 752 347 768 381
rect 802 347 818 381
rect -40 288 -6 347
rect 768 288 802 347
rect -40 -601 -6 -542
rect 768 -601 802 -542
rect -56 -635 -40 -601
rect -6 -635 10 -601
rect 752 -635 768 -601
rect 802 -635 818 -601
rect -140 -673 -106 -647
rect 868 -673 902 -647
rect -140 -707 -80 -673
rect 842 -707 902 -673
<< viali >>
rect -40 347 -6 381
rect 768 347 802 381
rect -40 -635 -6 -601
rect 768 -635 802 -601
<< metal1 >>
rect -52 381 6 387
rect -52 347 -40 381
rect -6 347 6 381
rect -52 341 6 347
rect 756 381 814 387
rect 756 347 768 381
rect 802 347 814 381
rect 756 341 814 347
rect -46 301 0 341
rect -46 299 88 301
rect 762 300 808 341
rect -60 101 -50 299
rect 4 101 88 299
rect 187 100 197 300
rect 249 100 259 300
rect 345 100 355 300
rect 407 100 417 300
rect 503 100 513 300
rect 565 100 575 300
rect 674 299 808 300
rect 674 100 758 299
rect 812 100 822 299
rect 97 -150 190 60
rect 302 13 460 59
rect 357 -15 403 13
rect 354 -21 406 -15
rect 354 -79 406 -73
rect 572 -150 664 59
rect 97 -199 348 -150
rect 35 -247 95 -241
rect 95 -307 191 -247
rect 35 -313 191 -307
rect 256 -312 348 -199
rect 414 -199 664 -150
rect 414 -312 506 -199
rect 667 -247 727 -241
rect 572 -307 667 -247
rect 572 -313 727 -307
rect -59 -554 -49 -354
rect 3 -554 86 -354
rect 187 -554 197 -354
rect 249 -554 259 -354
rect 344 -554 354 -356
rect 408 -554 418 -356
rect 503 -554 513 -354
rect 565 -554 575 -354
rect 674 -554 759 -354
rect 811 -554 821 -354
rect -46 -595 0 -554
rect 762 -595 808 -554
rect -52 -601 6 -595
rect -52 -635 -40 -601
rect -6 -635 6 -601
rect -52 -641 6 -635
rect 756 -601 814 -595
rect 756 -635 768 -601
rect 802 -635 814 -601
rect 756 -641 814 -635
<< via1 >>
rect -50 101 4 299
rect 197 100 249 300
rect 355 100 407 300
rect 513 100 565 300
rect 758 100 812 299
rect 354 -73 406 -21
rect 35 -307 95 -247
rect 667 -307 727 -247
rect -49 -554 3 -354
rect 197 -554 249 -354
rect 354 -554 408 -356
rect 513 -554 565 -354
rect 759 -554 811 -354
<< metal2 >>
rect 353 470 409 477
rect 351 468 411 470
rect 351 412 353 468
rect 409 412 411 468
rect -50 299 4 309
rect -284 212 -221 221
rect -284 -344 -221 149
rect -51 101 -50 299
rect -170 15 -161 75
rect -101 72 -92 75
rect -51 72 4 101
rect -101 17 4 72
rect 197 300 249 310
rect 351 300 411 412
rect 351 100 355 300
rect 407 100 411 300
rect 513 300 565 310
rect 565 100 566 300
rect -101 15 -92 17
rect 37 -46 93 -39
rect 35 -48 95 -46
rect 35 -104 37 -48
rect 93 -104 95 -48
rect 35 -247 95 -104
rect 197 -143 249 100
rect 355 90 407 100
rect 348 -46 354 -21
rect 406 -46 412 -21
rect 348 -73 350 -46
rect 410 -73 412 -46
rect 350 -115 410 -106
rect 513 -143 566 100
rect 758 299 812 309
rect 959 208 1019 217
rect 959 139 1019 148
rect 758 70 812 100
rect 864 75 924 84
rect 758 16 864 70
rect 924 16 926 70
rect 864 6 924 15
rect 669 -46 725 -39
rect 197 -189 566 -143
rect 29 -307 35 -247
rect 95 -307 101 -247
rect -284 -354 3 -344
rect -284 -407 -49 -354
rect -49 -564 3 -554
rect 197 -354 249 -189
rect 513 -306 566 -189
rect 667 -48 727 -46
rect 667 -104 669 -48
rect 725 -104 727 -48
rect 667 -247 727 -104
rect 354 -355 408 -346
rect 513 -354 565 -306
rect 661 -307 667 -247
rect 727 -307 733 -247
rect 967 -344 1010 139
rect 197 -564 249 -554
rect 351 -356 411 -355
rect 351 -554 354 -356
rect 408 -554 411 -356
rect 351 -703 411 -554
rect 513 -564 565 -554
rect 759 -354 1010 -344
rect 811 -407 1010 -354
rect 759 -564 811 -554
rect 344 -759 353 -703
rect 409 -759 418 -703
rect 351 -761 411 -759
<< via2 >>
rect 353 412 409 468
rect -284 149 -221 212
rect -161 15 -101 75
rect 37 -104 93 -48
rect 350 -73 354 -46
rect 354 -73 406 -46
rect 406 -73 410 -46
rect 350 -106 410 -73
rect 959 148 1019 208
rect 864 15 924 75
rect 669 -104 725 -48
rect 353 -759 409 -703
<< metal3 >>
rect -283 470 416 473
rect -283 468 1019 470
rect -283 412 353 468
rect 409 412 1019 468
rect -283 410 1019 412
rect -283 217 -220 410
rect 348 407 414 410
rect -289 212 -216 217
rect 959 213 1019 410
rect -289 149 -284 212
rect -221 149 -216 212
rect -289 144 -216 149
rect 954 208 1024 213
rect 954 148 959 208
rect 1019 148 1024 208
rect 954 143 1024 148
rect -166 75 -96 80
rect -166 15 -161 75
rect -101 15 -96 75
rect -166 10 -96 15
rect 859 75 929 80
rect 859 15 864 75
rect 924 15 929 75
rect 859 10 929 15
rect -161 -698 -101 10
rect 32 -46 98 -43
rect 345 -46 415 -41
rect 664 -46 730 -43
rect 32 -48 350 -46
rect 32 -104 37 -48
rect 93 -104 350 -48
rect 32 -106 350 -104
rect 410 -48 730 -46
rect 410 -104 669 -48
rect 725 -104 730 -48
rect 410 -106 730 -104
rect 32 -109 98 -106
rect 345 -111 415 -106
rect 664 -109 730 -106
rect -161 -701 414 -698
rect 864 -701 924 10
rect -161 -703 924 -701
rect -161 -758 353 -703
rect 348 -759 353 -758
rect 409 -759 924 -703
rect 348 -761 924 -759
rect 348 -764 414 -761
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729265743
transform 1 0 741 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729265743
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729265743
transform 1 0 21 0 1 -454
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729265743
transform 1 0 741 0 1 -454
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BH58Y6  sky130_fd_pr__pfet_01v8_BH58Y6_0
timestamp 1729265743
transform 1 0 381 0 1 -454
box -381 -200 381 200
use sky130_fd_pr__pfet_01v8_BH58Y6  sky130_fd_pr__pfet_01v8_BH58Y6_1
timestamp 1729265743
transform 1 0 381 0 1 200
box -381 -200 381 200
<< labels >>
flabel nsubdiffcont -121 279 -121 279 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel metal1 145 -159 145 -159 0 FreeSans 160 0 0 0 VIN
port 1 nsew
flabel metal2 -29 47 -29 47 0 FreeSans 160 0 0 0 D6
port 2 nsew
flabel metal2 226 73 226 73 0 FreeSans 160 0 0 0 D5
port 3 nsew
flabel metal3 450 -78 450 -78 0 FreeSans 160 0 0 0 VIP
port 4 nsew
flabel metal2 -254 14 -254 14 0 FreeSans 160 0 0 0 OUT
port 5 nsew
<< end >>
